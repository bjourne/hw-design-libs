library bjourne;
library ieee;
use ieee.numeric_std.all;

package types is
    type real_array2d_t is array(natural range<>) of real_vector;
end package;
