-- Copyright (C) 2023 Björn A. Lindqvist <bjourne@gmail.com>
library bjourne;
library ieee;
use bjourne.types.all;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity dct8x8 is
    port(
        clk, rstn : in std_logic;
        x : in real_array2d_t(0 to 7)(0 to 7);
        y : out real_array2d_t(0 to 7)(0 to 7)
    );
end dct8x8;

architecture rtl of dct8x8 is
    signal s1 : real_vector(0 to 63);
    signal s2 : real_vector(0 to 79);
    signal s3 : real_vector(0 to 87);
    signal s4 : real_vector(0 to 71);
    signal s5 : real_vector(0 to 63);
    signal s6 : real_vector(0 to 67);
    signal s7 : real_vector(0 to 69);
    signal s8 : real_vector(0 to 73);
    signal s9 : real_vector(0 to 79);
    signal s10 : real_vector(0 to 73);
    signal s11 : real_vector(0 to 65);
    signal s12 : real_vector(0 to 63);
    signal s13 : real_vector(0 to 63);
    signal s14 : real_vector(0 to 63);
begin
    y <= (
        (s14(4), s14(5), s14(6), s14(7), s14(8), s14(9), s14(10), s14(11)),
        (s14(12), s14(0), s14(13), s14(14), s14(15), s14(16), s14(17), s14(1)),
        (s14(18), s14(19), s14(20), s14(21), s14(22), s14(23), s14(24), s14(25)),
        (s14(26), s14(27), s14(28), s14(29), s14(30), s14(31), s14(32), s14(33)),
        (s14(34), s14(35), s14(36), s14(37), s14(38), s14(39), s14(40), s14(41)),
        (s14(42), s14(43), s14(44), s14(45), s14(46), s14(47), s14(48), s14(49)),
        (s14(50), s14(51), s14(52), s14(53), s14(54), s14(55), s14(56), s14(57)),
        (s14(58), s14(2), s14(59), s14(60), s14(61), s14(62), s14(63), s14(3))
    );
    process (clk)
    begin
        if rising_edge(clk) then
            if rstn = '0' then
                s1 <= (others => 0.0);
                s2 <= (others => 0.0);
                s3 <= (others => 0.0);
                s4 <= (others => 0.0);
                s5 <= (others => 0.0);
                s6 <= (others => 0.0);
                s7 <= (others => 0.0);
                s8 <= (others => 0.0);
                s9 <= (others => 0.0);
                s10 <= (others => 0.0);
                s11 <= (others => 0.0);
                s12 <= (others => 0.0);
                s13 <= (others => 0.0);
                s14 <= (others => 0.0);
            else
                s1(0)  <= x(0)(0) + x(0)(7);
                s1(1)  <= x(0)(3) + x(0)(4);
                s1(2)  <= x(0)(1) + x(0)(6);
                s1(3)  <= x(0)(2) + x(0)(5);
                s1(4)  <= x(7)(0) + x(7)(7);
                s1(5)  <= x(7)(3) + x(7)(4);
                s1(6)  <= x(7)(1) + x(7)(6);
                s1(7)  <= x(7)(2) + x(7)(5);
                s1(8)  <= x(3)(0) + x(3)(7);
                s1(9)  <= x(3)(3) + x(3)(4);
                s1(10) <= x(3)(1) + x(3)(6);
                s1(11) <= x(3)(2) + x(3)(5);
                s1(12) <= x(4)(0) + x(4)(7);
                s1(13) <= x(4)(3) + x(4)(4);
                s1(14) <= x(4)(1) + x(4)(6);
                s1(15) <= x(4)(2) + x(4)(5);
                s1(16) <= x(1)(0) + x(1)(7);
                s1(17) <= x(1)(3) + x(1)(4);
                s1(18) <= x(1)(1) + x(1)(6);
                s1(19) <= x(1)(2) + x(1)(5);
                s1(20) <= x(6)(0) + x(6)(7);
                s1(21) <= x(6)(3) + x(6)(4);
                s1(22) <= x(6)(1) + x(6)(6);
                s1(23) <= x(6)(2) + x(6)(5);
                s1(24) <= x(2)(0) + x(2)(7);
                s1(25) <= x(2)(3) + x(2)(4);
                s1(26) <= x(2)(1) + x(2)(6);
                s1(27) <= x(2)(2) + x(2)(5);
                s1(28) <= x(5)(0) + x(5)(7);
                s1(29) <= x(5)(3) + x(5)(4);
                s1(30) <= x(5)(1) + x(5)(6);
                s1(31) <= x(5)(2) + x(5)(5);
                s1(32) <= x(0)(3) - x(0)(4);
                s1(33) <= x(0)(0) - x(0)(7);
                s1(34) <= x(0)(1) - x(0)(6);
                s1(35) <= x(0)(2) - x(0)(5);
                s1(36) <= x(7)(3) - x(7)(4);
                s1(37) <= x(7)(0) - x(7)(7);
                s1(38) <= x(7)(1) - x(7)(6);
                s1(39) <= x(7)(2) - x(7)(5);
                s1(40) <= x(3)(3) - x(3)(4);
                s1(41) <= x(3)(0) - x(3)(7);
                s1(42) <= x(3)(1) - x(3)(6);
                s1(43) <= x(3)(2) - x(3)(5);
                s1(44) <= x(4)(3) - x(4)(4);
                s1(45) <= x(4)(0) - x(4)(7);
                s1(46) <= x(4)(1) - x(4)(6);
                s1(47) <= x(4)(2) - x(4)(5);
                s1(48) <= x(1)(3) - x(1)(4);
                s1(49) <= x(1)(0) - x(1)(7);
                s1(50) <= x(1)(1) - x(1)(6);
                s1(51) <= x(1)(2) - x(1)(5);
                s1(52) <= x(6)(3) - x(6)(4);
                s1(53) <= x(6)(0) - x(6)(7);
                s1(54) <= x(6)(1) - x(6)(6);
                s1(55) <= x(6)(2) - x(6)(5);
                s1(56) <= x(2)(3) - x(2)(4);
                s1(57) <= x(2)(0) - x(2)(7);
                s1(58) <= x(2)(1) - x(2)(6);
                s1(59) <= x(2)(2) - x(2)(5);
                s1(60) <= x(5)(3) - x(5)(4);
                s1(61) <= x(5)(0) - x(5)(7);
                s1(62) <= x(5)(1) - x(5)(6);
                s1(63) <= x(5)(2) - x(5)(5);
                s2(0)  <= s1(0) + s1(1);
                s2(1)  <= s1(2) + s1(3);
                s2(2)  <= s1(4) + s1(5);
                s2(3)  <= s1(6) + s1(7);
                s2(4)  <= s1(8) + s1(9);
                s2(5)  <= s1(10) + s1(11);
                s2(6)  <= s1(12) + s1(13);
                s2(7)  <= s1(14) + s1(15);
                s2(8)  <= s1(16) + s1(17);
                s2(9)  <= s1(18) + s1(19);
                s2(10) <= s1(20) + s1(21);
                s2(11) <= s1(22) + s1(23);
                s2(12) <= s1(24) + s1(25);
                s2(13) <= s1(26) + s1(27);
                s2(14) <= s1(28) + s1(29);
                s2(15) <= s1(30) + s1(31);
                s2(16) <= -1.38703984532 * s1(32);
                s2(17) <= s1(32) + s1(33);
                s2(18) <= -0.78569495838 * s1(34);
                s2(19) <= s1(35) + s1(34);
                s2(20) <= -0.27589937928 * s1(33);
                s2(21) <= -1.17587560241 * s1(35);
                s2(22) <= -1.38703984532 * s1(36);
                s2(23) <= s1(36) + s1(37);
                s2(24) <= -0.78569495838 * s1(38);
                s2(25) <= s1(39) + s1(38);
                s2(26) <= -0.27589937928 * s1(37);
                s2(27) <= -1.17587560241 * s1(39);
                s2(28) <= -1.38703984532 * s1(40);
                s2(29) <= s1(40) + s1(41);
                s2(30) <= -0.78569495838 * s1(42);
                s2(31) <= s1(43) + s1(42);
                s2(32) <= -0.27589937928 * s1(41);
                s2(33) <= -1.17587560241 * s1(43);
                s2(34) <= -1.38703984532 * s1(44);
                s2(35) <= s1(44) + s1(45);
                s2(36) <= -0.78569495838 * s1(46);
                s2(37) <= s1(47) + s1(46);
                s2(38) <= -0.27589937928 * s1(45);
                s2(39) <= -1.17587560241 * s1(47);
                s2(40) <= -1.38703984532 * s1(48);
                s2(41) <= s1(48) + s1(49);
                s2(42) <= -0.78569495838 * s1(50);
                s2(43) <= s1(51) + s1(50);
                s2(44) <= -0.27589937928 * s1(49);
                s2(45) <= -1.17587560241 * s1(51);
                s2(46) <= -1.38703984532 * s1(52);
                s2(47) <= s1(52) + s1(53);
                s2(48) <= -0.78569495838 * s1(54);
                s2(49) <= s1(55) + s1(54);
                s2(50) <= -0.27589937928 * s1(53);
                s2(51) <= -1.17587560241 * s1(55);
                s2(52) <= -1.38703984532 * s1(56);
                s2(53) <= s1(56) + s1(57);
                s2(54) <= -0.78569495838 * s1(58);
                s2(55) <= s1(59) + s1(58);
                s2(56) <= -0.27589937928 * s1(57);
                s2(57) <= -1.17587560241 * s1(59);
                s2(58) <= -1.38703984532 * s1(60);
                s2(59) <= s1(60) + s1(61);
                s2(60) <= -0.78569495838 * s1(62);
                s2(61) <= s1(63) + s1(62);
                s2(62) <= -0.27589937928 * s1(61);
                s2(63) <= -1.17587560241 * s1(63);
                s2(64) <= s1(0) - s1(1);
                s2(65) <= s1(2) - s1(3);
                s2(66) <= s1(4) - s1(5);
                s2(67) <= s1(6) - s1(7);
                s2(68) <= s1(8) - s1(9);
                s2(69) <= s1(10) - s1(11);
                s2(70) <= s1(12) - s1(13);
                s2(71) <= s1(14) - s1(15);
                s2(72) <= s1(16) - s1(17);
                s2(73) <= s1(18) - s1(19);
                s2(74) <= s1(20) - s1(21);
                s2(75) <= s1(22) - s1(23);
                s2(76) <= s1(24) - s1(25);
                s2(77) <= s1(26) - s1(27);
                s2(78) <= s1(28) - s1(29);
                s2(79) <= s1(30) - s1(31);
                s3(0)  <= s2(0) + s2(1);
                s3(1)  <= s2(2) + s2(3);
                s3(2)  <= s2(4) + s2(5);
                s3(3)  <= s2(6) + s2(7);
                s3(4)  <= s2(8) + s2(9);
                s3(5)  <= s2(10) + s2(11);
                s3(6)  <= s2(12) + s2(13);
                s3(7)  <= s2(14) + s2(15);
                s3(8)  <= 0.8314696123 * s2(17);
                s3(9)  <= 0.9807852804 * s2(19);
                s3(10) <= 0.8314696123 * s2(23);
                s3(11) <= 0.9807852804 * s2(25);
                s3(12) <= 0.8314696123 * s2(29);
                s3(13) <= 0.9807852804 * s2(31);
                s3(14) <= 0.8314696123 * s2(35);
                s3(15) <= 0.9807852804 * s2(37);
                s3(16) <= 0.8314696123 * s2(41);
                s3(17) <= 0.9807852804 * s2(43);
                s3(18) <= 0.8314696123 * s2(47);
                s3(19) <= 0.9807852804 * s2(49);
                s3(20) <= 0.8314696123 * s2(53);
                s3(21) <= 0.9807852804 * s2(55);
                s3(22) <= 0.8314696123 * s2(59);
                s3(23) <= 0.9807852804 * s2(61);
                s3(24) <= 0.76536686473 * s2(64);
                s3(25) <= s2(65) + s2(64);
                s3(26) <= 0.76536686473 * s2(66);
                s3(27) <= s2(67) + s2(66);
                s3(28) <= 0.76536686473 * s2(68);
                s3(29) <= s2(69) + s2(68);
                s3(30) <= 0.76536686473 * s2(70);
                s3(31) <= s2(71) + s2(70);
                s3(32) <= 0.76536686473 * s2(72);
                s3(33) <= s2(73) + s2(72);
                s3(34) <= 0.76536686473 * s2(74);
                s3(35) <= s2(75) + s2(74);
                s3(36) <= 0.76536686473 * s2(76);
                s3(37) <= s2(77) + s2(76);
                s3(38) <= 0.76536686473 * s2(78);
                s3(39) <= s2(79) + s2(78);
                s3(40) <= s2(0) - s2(1);
                s3(41) <= s2(2) - s2(3);
                s3(42) <= s2(4) - s2(5);
                s3(43) <= s2(6) - s2(7);
                s3(44) <= s2(8) - s2(9);
                s3(45) <= s2(10) - s2(11);
                s3(46) <= s2(12) - s2(13);
                s3(47) <= s2(14) - s2(15);
                s3(48) <= -1.84775906502 * s2(65);
                s3(49) <= -1.84775906502 * s2(67);
                s3(50) <= -1.84775906502 * s2(69);
                s3(51) <= -1.84775906502 * s2(71);
                s3(52) <= -1.84775906502 * s2(73);
                s3(53) <= -1.84775906502 * s2(75);
                s3(54) <= -1.84775906502 * s2(77);
                s3(55) <= -1.84775906502 * s2(79);
                s3(56) <= s2(16);
                s3(57) <= s2(18);
                s3(58) <= s2(20);
                s3(59) <= s2(21);
                s3(60) <= s2(22);
                s3(61) <= s2(24);
                s3(62) <= s2(26);
                s3(63) <= s2(27);
                s3(64) <= s2(28);
                s3(65) <= s2(30);
                s3(66) <= s2(32);
                s3(67) <= s2(33);
                s3(68) <= s2(34);
                s3(69) <= s2(36);
                s3(70) <= s2(38);
                s3(71) <= s2(39);
                s3(72) <= s2(40);
                s3(73) <= s2(42);
                s3(74) <= s2(44);
                s3(75) <= s2(45);
                s3(76) <= s2(46);
                s3(77) <= s2(48);
                s3(78) <= s2(50);
                s3(79) <= s2(51);
                s3(80) <= s2(52);
                s3(81) <= s2(54);
                s3(82) <= s2(56);
                s3(83) <= s2(57);
                s3(84) <= s2(58);
                s3(85) <= s2(60);
                s3(86) <= s2(62);
                s3(87) <= s2(63);
                s4(0)  <= 0.35355339059 * s3(0);
                s4(1)  <= 0.35355339059 * s3(1);
                s4(2)  <= 0.35355339059 * s3(2);
                s4(3)  <= 0.35355339059 * s3(3);
                s4(4)  <= 0.35355339059 * s3(4);
                s4(5)  <= 0.35355339059 * s3(5);
                s4(6)  <= 0.35355339059 * s3(6);
                s4(7)  <= 0.35355339059 * s3(7);
                s4(8)  <= s3(56) + s3(8);
                s4(9)  <= s3(57) + s3(9);
                s4(10) <= s3(58) + s3(8);
                s4(11) <= s3(59) + s3(9);
                s4(12) <= s3(60) + s3(10);
                s4(13) <= s3(61) + s3(11);
                s4(14) <= s3(62) + s3(10);
                s4(15) <= s3(63) + s3(11);
                s4(16) <= s3(64) + s3(12);
                s4(17) <= s3(65) + s3(13);
                s4(18) <= s3(66) + s3(12);
                s4(19) <= s3(67) + s3(13);
                s4(20) <= s3(68) + s3(14);
                s4(21) <= s3(69) + s3(15);
                s4(22) <= s3(70) + s3(14);
                s4(23) <= s3(71) + s3(15);
                s4(24) <= s3(72) + s3(16);
                s4(25) <= s3(73) + s3(17);
                s4(26) <= s3(74) + s3(16);
                s4(27) <= s3(75) + s3(17);
                s4(28) <= s3(76) + s3(18);
                s4(29) <= s3(77) + s3(19);
                s4(30) <= s3(78) + s3(18);
                s4(31) <= s3(79) + s3(19);
                s4(32) <= s3(80) + s3(20);
                s4(33) <= s3(81) + s3(21);
                s4(34) <= s3(82) + s3(20);
                s4(35) <= s3(83) + s3(21);
                s4(36) <= s3(84) + s3(22);
                s4(37) <= s3(85) + s3(23);
                s4(38) <= s3(86) + s3(22);
                s4(39) <= s3(87) + s3(23);
                s4(40) <= 0.54119610014 * s3(25);
                s4(41) <= 0.54119610014 * s3(27);
                s4(42) <= 0.54119610014 * s3(29);
                s4(43) <= 0.54119610014 * s3(31);
                s4(44) <= 0.54119610014 * s3(33);
                s4(45) <= 0.54119610014 * s3(35);
                s4(46) <= 0.54119610014 * s3(37);
                s4(47) <= 0.54119610014 * s3(39);
                s4(48) <= 0.35355339059 * s3(40);
                s4(49) <= 0.35355339059 * s3(41);
                s4(50) <= 0.35355339059 * s3(42);
                s4(51) <= 0.35355339059 * s3(43);
                s4(52) <= 0.35355339059 * s3(44);
                s4(53) <= 0.35355339059 * s3(45);
                s4(54) <= 0.35355339059 * s3(46);
                s4(55) <= 0.35355339059 * s3(47);
                s4(56) <= s3(24);
                s4(57) <= s3(26);
                s4(58) <= s3(28);
                s4(59) <= s3(30);
                s4(60) <= s3(32);
                s4(61) <= s3(34);
                s4(62) <= s3(36);
                s4(63) <= s3(38);
                s4(64) <= s3(48);
                s4(65) <= s3(49);
                s4(66) <= s3(50);
                s4(67) <= s3(51);
                s4(68) <= s3(52);
                s4(69) <= s3(53);
                s4(70) <= s3(54);
                s4(71) <= s3(55);
                s5(0)  <= s4(0) + s4(1);
                s5(1)  <= s4(2) + s4(3);
                s5(2)  <= s4(4) + s4(5);
                s5(3)  <= s4(6) + s4(7);
                s5(4)  <= s4(8) + s4(9);
                s5(5)  <= s4(10) + s4(11);
                s5(6)  <= s4(12) + s4(13);
                s5(7)  <= s4(14) + s4(15);
                s5(8)  <= s4(16) + s4(17);
                s5(9)  <= s4(18) + s4(19);
                s5(10) <= s4(20) + s4(21);
                s5(11) <= s4(22) + s4(23);
                s5(12) <= s4(24) + s4(25);
                s5(13) <= s4(26) + s4(27);
                s5(14) <= s4(28) + s4(29);
                s5(15) <= s4(30) + s4(31);
                s5(16) <= s4(32) + s4(33);
                s5(17) <= s4(34) + s4(35);
                s5(18) <= s4(36) + s4(37);
                s5(19) <= s4(38) + s4(39);
                s5(20) <= s4(56) + s4(40);
                s5(21) <= s4(57) + s4(41);
                s5(22) <= s4(58) + s4(42);
                s5(23) <= s4(59) + s4(43);
                s5(24) <= s4(60) + s4(44);
                s5(25) <= s4(61) + s4(45);
                s5(26) <= s4(62) + s4(46);
                s5(27) <= s4(63) + s4(47);
                s5(28) <= s4(8) - s4(9);
                s5(29) <= s4(12) - s4(13);
                s5(30) <= s4(16) - s4(17);
                s5(31) <= s4(20) - s4(21);
                s5(32) <= s4(24) - s4(25);
                s5(33) <= s4(28) - s4(29);
                s5(34) <= s4(32) - s4(33);
                s5(35) <= s4(36) - s4(37);
                s5(36) <= s4(48) + s4(49);
                s5(37) <= s4(50) + s4(51);
                s5(38) <= s4(52) + s4(53);
                s5(39) <= s4(54) + s4(55);
                s5(40) <= s4(10) - s4(11);
                s5(41) <= s4(14) - s4(15);
                s5(42) <= s4(18) - s4(19);
                s5(43) <= s4(22) - s4(23);
                s5(44) <= s4(26) - s4(27);
                s5(45) <= s4(30) - s4(31);
                s5(46) <= s4(34) - s4(35);
                s5(47) <= s4(38) - s4(39);
                s5(48) <= s4(64) + s4(40);
                s5(49) <= s4(65) + s4(41);
                s5(50) <= s4(66) + s4(42);
                s5(51) <= s4(67) + s4(43);
                s5(52) <= s4(68) + s4(44);
                s5(53) <= s4(69) + s4(45);
                s5(54) <= s4(70) + s4(46);
                s5(55) <= s4(71) + s4(47);
                s5(56) <= s4(2) - s4(3);
                s5(57) <= s4(0) - s4(1);
                s5(58) <= s4(4) - s4(5);
                s5(59) <= s4(6) - s4(7);
                s5(60) <= s4(50) - s4(51);
                s5(61) <= s4(48) - s4(49);
                s5(62) <= s4(52) - s4(53);
                s5(63) <= s4(54) - s4(55);
                s6(0)  <= s5(0) + s5(1);
                s6(1)  <= s5(2) + s5(3);
                s6(2)  <= s5(4) + s5(5);
                s6(3)  <= s5(6) + s5(7);
                s6(4)  <= s5(8) + s5(9);
                s6(5)  <= s5(10) + s5(11);
                s6(6)  <= s5(12) + s5(13);
                s6(7)  <= s5(14) + s5(15);
                s6(8)  <= s5(16) + s5(17);
                s6(9)  <= s5(18) + s5(19);
                s6(10) <= 0.35355339059 * s5(20);
                s6(11) <= 0.35355339059 * s5(21);
                s6(12) <= 0.35355339059 * s5(22);
                s6(13) <= 0.35355339059 * s5(23);
                s6(14) <= 0.35355339059 * s5(24);
                s6(15) <= 0.35355339059 * s5(25);
                s6(16) <= 0.35355339059 * s5(26);
                s6(17) <= 0.35355339059 * s5(27);
                s6(18) <= 0.5 * s5(28);
                s6(19) <= 0.5 * s5(29);
                s6(20) <= 0.5 * s5(30);
                s6(21) <= 0.5 * s5(31);
                s6(22) <= 0.5 * s5(32);
                s6(23) <= 0.5 * s5(33);
                s6(24) <= 0.5 * s5(34);
                s6(25) <= 0.5 * s5(35);
                s6(26) <= s5(36) + s5(37);
                s6(27) <= s5(38) + s5(39);
                s6(28) <= 0.5 * s5(40);
                s6(29) <= 0.5 * s5(41);
                s6(30) <= 0.5 * s5(42);
                s6(31) <= 0.5 * s5(43);
                s6(32) <= 0.5 * s5(44);
                s6(33) <= 0.5 * s5(45);
                s6(34) <= 0.5 * s5(46);
                s6(35) <= 0.5 * s5(47);
                s6(36) <= 0.35355339059 * s5(48);
                s6(37) <= 0.35355339059 * s5(49);
                s6(38) <= 0.35355339059 * s5(50);
                s6(39) <= 0.35355339059 * s5(51);
                s6(40) <= 0.35355339059 * s5(52);
                s6(41) <= 0.35355339059 * s5(53);
                s6(42) <= 0.35355339059 * s5(54);
                s6(43) <= 0.35355339059 * s5(55);
                s6(44) <= s5(4) - s5(5);
                s6(45) <= s5(6) - s5(7);
                s6(46) <= s5(8) - s5(9);
                s6(47) <= s5(10) - s5(11);
                s6(48) <= s5(12) - s5(13);
                s6(49) <= s5(14) - s5(15);
                s6(50) <= s5(16) - s5(17);
                s6(51) <= s5(18) - s5(19);
                s6(52) <= -1.38703984532 * s5(56);
                s6(53) <= s5(56) + s5(57);
                s6(54) <= -0.78569495838 * s5(58);
                s6(55) <= s5(59) + s5(58);
                s6(56) <= -0.27589937928 * s5(57);
                s6(57) <= -1.17587560241 * s5(59);
                s6(58) <= -1.38703984532 * s5(60);
                s6(59) <= s5(60) + s5(61);
                s6(60) <= -0.78569495838 * s5(62);
                s6(61) <= s5(63) + s5(62);
                s6(62) <= -0.27589937928 * s5(61);
                s6(63) <= -1.17587560241 * s5(63);
                s6(64) <= s5(0) - s5(1);
                s6(65) <= s5(2) - s5(3);
                s6(66) <= s5(36) - s5(37);
                s6(67) <= s5(38) - s5(39);
                s7(0)  <= s6(0) + s6(1);
                s7(1)  <= 0.35355339059 * s6(2);
                s7(2)  <= 0.35355339059 * s6(3);
                s7(3)  <= 0.35355339059 * s6(4);
                s7(4)  <= 0.35355339059 * s6(5);
                s7(5)  <= 0.35355339059 * s6(6);
                s7(6)  <= 0.35355339059 * s6(7);
                s7(7)  <= 0.35355339059 * s6(8);
                s7(8)  <= 0.35355339059 * s6(9);
                s7(9)  <= s6(10) + s6(11);
                s7(10) <= s6(12) + s6(13);
                s7(11) <= s6(14) + s6(15);
                s7(12) <= s6(16) + s6(17);
                s7(13) <= s6(18) + s6(19);
                s7(14) <= s6(20) + s6(21);
                s7(15) <= s6(22) + s6(23);
                s7(16) <= s6(24) + s6(25);
                s7(17) <= s6(26) + s6(27);
                s7(18) <= s6(28) + s6(29);
                s7(19) <= s6(30) + s6(31);
                s7(20) <= s6(32) + s6(33);
                s7(21) <= s6(34) + s6(35);
                s7(22) <= s6(36) + s6(37);
                s7(23) <= s6(38) + s6(39);
                s7(24) <= s6(40) + s6(41);
                s7(25) <= s6(42) + s6(43);
                s7(26) <= 0.35355339059 * s6(44);
                s7(27) <= 0.35355339059 * s6(45);
                s7(28) <= 0.35355339059 * s6(46);
                s7(29) <= 0.35355339059 * s6(47);
                s7(30) <= 0.35355339059 * s6(48);
                s7(31) <= 0.35355339059 * s6(49);
                s7(32) <= 0.35355339059 * s6(50);
                s7(33) <= 0.35355339059 * s6(51);
                s7(34) <= 0.8314696123 * s6(53);
                s7(35) <= 0.9807852804 * s6(55);
                s7(36) <= s6(12) - s6(13);
                s7(37) <= s6(10) - s6(11);
                s7(38) <= s6(14) - s6(15);
                s7(39) <= s6(16) - s6(17);
                s7(40) <= s6(20) - s6(21);
                s7(41) <= s6(18) - s6(19);
                s7(42) <= s6(22) - s6(23);
                s7(43) <= s6(24) - s6(25);
                s7(44) <= 0.8314696123 * s6(59);
                s7(45) <= 0.9807852804 * s6(61);
                s7(46) <= s6(30) - s6(31);
                s7(47) <= s6(28) - s6(29);
                s7(48) <= s6(32) - s6(33);
                s7(49) <= s6(34) - s6(35);
                s7(50) <= s6(38) - s6(39);
                s7(51) <= s6(36) - s6(37);
                s7(52) <= s6(40) - s6(41);
                s7(53) <= s6(42) - s6(43);
                s7(54) <= 0.76536686473 * s6(64);
                s7(55) <= s6(65) + s6(64);
                s7(56) <= 0.76536686473 * s6(66);
                s7(57) <= s6(67) + s6(66);
                s7(58) <= s6(0) - s6(1);
                s7(59) <= s6(26) - s6(27);
                s7(60) <= -1.84775906502 * s6(65);
                s7(61) <= -1.84775906502 * s6(67);
                s7(62) <= s6(52);
                s7(63) <= s6(54);
                s7(64) <= s6(56);
                s7(65) <= s6(57);
                s7(66) <= s6(58);
                s7(67) <= s6(60);
                s7(68) <= s6(62);
                s7(69) <= s6(63);
                s8(0)  <= 0.35355339059 * s7(0);
                s8(1)  <= s7(1) + s7(2);
                s8(2)  <= s7(3) + s7(4);
                s8(3)  <= s7(5) + s7(6);
                s8(4)  <= s7(7) + s7(8);
                s8(5)  <= s7(9) + s7(10);
                s8(6)  <= s7(11) + s7(12);
                s8(7)  <= s7(13) + s7(14);
                s8(8)  <= s7(15) + s7(16);
                s8(9)  <= 0.35355339059 * s7(17);
                s8(10) <= s7(18) + s7(19);
                s8(11) <= s7(20) + s7(21);
                s8(12) <= s7(22) + s7(23);
                s8(13) <= s7(24) + s7(25);
                s8(14) <= s7(26) + s7(27);
                s8(15) <= s7(28) + s7(29);
                s8(16) <= s7(30) + s7(31);
                s8(17) <= s7(32) + s7(33);
                s8(18) <= s7(62) + s7(34);
                s8(19) <= s7(63) + s7(35);
                s8(20) <= s7(64) + s7(34);
                s8(21) <= s7(65) + s7(35);
                s8(22) <= s7(3) - s7(4);
                s8(23) <= s7(1) - s7(2);
                s8(24) <= s7(5) - s7(6);
                s8(25) <= s7(7) - s7(8);
                s8(26) <= -1.38703984532 * s7(36);
                s8(27) <= s7(36) + s7(37);
                s8(28) <= -0.78569495838 * s7(38);
                s8(29) <= s7(39) + s7(38);
                s8(30) <= -0.27589937928 * s7(37);
                s8(31) <= -1.17587560241 * s7(39);
                s8(32) <= -1.38703984532 * s7(40);
                s8(33) <= s7(40) + s7(41);
                s8(34) <= -0.78569495838 * s7(42);
                s8(35) <= s7(43) + s7(42);
                s8(36) <= -0.27589937928 * s7(41);
                s8(37) <= -1.17587560241 * s7(43);
                s8(38) <= s7(66) + s7(44);
                s8(39) <= s7(67) + s7(45);
                s8(40) <= s7(68) + s7(44);
                s8(41) <= s7(69) + s7(45);
                s8(42) <= -1.38703984532 * s7(46);
                s8(43) <= s7(46) + s7(47);
                s8(44) <= -0.78569495838 * s7(48);
                s8(45) <= s7(49) + s7(48);
                s8(46) <= -0.27589937928 * s7(47);
                s8(47) <= -1.17587560241 * s7(49);
                s8(48) <= -1.38703984532 * s7(50);
                s8(49) <= s7(50) + s7(51);
                s8(50) <= -0.78569495838 * s7(52);
                s8(51) <= s7(53) + s7(52);
                s8(52) <= -0.27589937928 * s7(51);
                s8(53) <= -1.17587560241 * s7(53);
                s8(54) <= s7(28) - s7(29);
                s8(55) <= s7(26) - s7(27);
                s8(56) <= s7(30) - s7(31);
                s8(57) <= s7(32) - s7(33);
                s8(58) <= 0.54119610014 * s7(55);
                s8(59) <= s7(9) - s7(10);
                s8(60) <= s7(11) - s7(12);
                s8(61) <= s7(13) - s7(14);
                s8(62) <= s7(15) - s7(16);
                s8(63) <= 0.54119610014 * s7(57);
                s8(64) <= s7(18) - s7(19);
                s8(65) <= s7(20) - s7(21);
                s8(66) <= s7(22) - s7(23);
                s8(67) <= s7(24) - s7(25);
                s8(68) <= 0.35355339059 * s7(58);
                s8(69) <= 0.35355339059 * s7(59);
                s8(70) <= s7(54);
                s8(71) <= s7(56);
                s8(72) <= s7(60);
                s8(73) <= s7(61);
                s9(0)  <= s8(1) + s8(2);
                s9(1)  <= s8(3) + s8(4);
                s9(2)  <= s8(5) + s8(6);
                s9(3)  <= s8(7) + s8(8);
                s9(4)  <= s8(10) + s8(11);
                s9(5)  <= s8(12) + s8(13);
                s9(6)  <= s8(14) + s8(15);
                s9(7)  <= s8(16) + s8(17);
                s9(8)  <= s8(18) + s8(19);
                s9(9)  <= s8(20) + s8(21);
                s9(10) <= -1.38703984532 * s8(22);
                s9(11) <= s8(22) + s8(23);
                s9(12) <= -0.78569495838 * s8(24);
                s9(13) <= s8(25) + s8(24);
                s9(14) <= -0.27589937928 * s8(23);
                s9(15) <= -1.17587560241 * s8(25);
                s9(16) <= 0.8314696123 * s8(27);
                s9(17) <= 0.9807852804 * s8(29);
                s9(18) <= 0.8314696123 * s8(33);
                s9(19) <= 0.9807852804 * s8(35);
                s9(20) <= s8(38) + s8(39);
                s9(21) <= s8(40) + s8(41);
                s9(22) <= 0.8314696123 * s8(43);
                s9(23) <= 0.9807852804 * s8(45);
                s9(24) <= 0.8314696123 * s8(49);
                s9(25) <= 0.9807852804 * s8(51);
                s9(26) <= -1.38703984532 * s8(54);
                s9(27) <= s8(54) + s8(55);
                s9(28) <= -0.78569495838 * s8(56);
                s9(29) <= s8(57) + s8(56);
                s9(30) <= -0.27589937928 * s8(55);
                s9(31) <= -1.17587560241 * s8(57);
                s9(32) <= s8(70) + s8(58);
                s9(33) <= s8(1) - s8(2);
                s9(34) <= s8(3) - s8(4);
                s9(35) <= 0.76536686473 * s8(59);
                s9(36) <= s8(60) + s8(59);
                s9(37) <= 0.76536686473 * s8(61);
                s9(38) <= s8(62) + s8(61);
                s9(39) <= s8(71) + s8(63);
                s9(40) <= 0.76536686473 * s8(64);
                s9(41) <= s8(65) + s8(64);
                s9(42) <= 0.76536686473 * s8(66);
                s9(43) <= s8(67) + s8(66);
                s9(44) <= s8(14) - s8(15);
                s9(45) <= s8(16) - s8(17);
                s9(46) <= s8(18) - s8(19);
                s9(47) <= s8(38) - s8(39);
                s9(48) <= s8(5) - s8(6);
                s9(49) <= s8(7) - s8(8);
                s9(50) <= s8(10) - s8(11);
                s9(51) <= s8(12) - s8(13);
                s9(52) <= s8(20) - s8(21);
                s9(53) <= s8(40) - s8(41);
                s9(54) <= s8(72) + s8(58);
                s9(55) <= -1.84775906502 * s8(60);
                s9(56) <= -1.84775906502 * s8(62);
                s9(57) <= s8(73) + s8(63);
                s9(58) <= -1.84775906502 * s8(65);
                s9(59) <= -1.84775906502 * s8(67);
                s9(60) <= s8(0);
                s9(61) <= s8(9);
                s9(62) <= s8(26);
                s9(63) <= s8(28);
                s9(64) <= s8(30);
                s9(65) <= s8(31);
                s9(66) <= s8(32);
                s9(67) <= s8(34);
                s9(68) <= s8(36);
                s9(69) <= s8(37);
                s9(70) <= s8(42);
                s9(71) <= s8(44);
                s9(72) <= s8(46);
                s9(73) <= s8(47);
                s9(74) <= s8(48);
                s9(75) <= s8(50);
                s9(76) <= s8(52);
                s9(77) <= s8(53);
                s9(78) <= s8(68);
                s9(79) <= s8(69);
                s10(0) <= s9(0) + s9(1);
                s10(1) <= 0.35355339059 * s9(2);
                s10(2) <= 0.35355339059 * s9(3);
                s10(3) <= 0.35355339059 * s9(4);
                s10(4) <= 0.35355339059 * s9(5);
                s10(5) <= s9(6) + s9(7);
                s10(6) <= s9(8) + s9(9);
                s10(7) <= 0.8314696123 * s9(11);
                s10(8) <= 0.9807852804 * s9(13);
                s10(9) <= s9(62) + s9(16);
                s10(10) <= s9(63) + s9(17);
                s10(11) <= s9(64) + s9(16);
                s10(12) <= s9(65) + s9(17);
                s10(13) <= s9(66) + s9(18);
                s10(14) <= s9(67) + s9(19);
                s10(15) <= s9(68) + s9(18);
                s10(16) <= s9(69) + s9(19);
                s10(17) <= s9(20) + s9(21);
                s10(18) <= s9(70) + s9(22);
                s10(19) <= s9(71) + s9(23);
                s10(20) <= s9(72) + s9(22);
                s10(21) <= s9(73) + s9(23);
                s10(22) <= s9(74) + s9(24);
                s10(23) <= s9(75) + s9(25);
                s10(24) <= s9(76) + s9(24);
                s10(25) <= s9(77) + s9(25);
                s10(26) <= 0.8314696123 * s9(27);
                s10(27) <= 0.9807852804 * s9(29);
                s10(28) <= 0.35355339059 * s9(32);
                s10(29) <= 0.76536686473 * s9(33);
                s10(30) <= s9(34) + s9(33);
                s10(31) <= 0.54119610014 * s9(36);
                s10(32) <= 0.54119610014 * s9(38);
                s10(33) <= 0.35355339059 * s9(39);
                s10(34) <= 0.54119610014 * s9(41);
                s10(35) <= 0.54119610014 * s9(43);
                s10(36) <= 0.76536686473 * s9(44);
                s10(37) <= s9(45) + s9(44);
                s10(38) <= 0.5 * s9(46);
                s10(39) <= 0.5 * s9(47);
                s10(40) <= s9(0) - s9(1);
                s10(41) <= 0.35355339059 * s9(48);
                s10(42) <= 0.35355339059 * s9(49);
                s10(43) <= 0.35355339059 * s9(50);
                s10(44) <= 0.35355339059 * s9(51);
                s10(45) <= s9(6) - s9(7);
                s10(46) <= 0.5 * s9(52);
                s10(47) <= 0.5 * s9(53);
                s10(48) <= 0.35355339059 * s9(54);
                s10(49) <= -1.84775906502 * s9(34);
                s10(50) <= 0.35355339059 * s9(57);
                s10(51) <= -1.84775906502 * s9(45);
                s10(52) <= s9(8) - s9(9);
                s10(53) <= s9(20) - s9(21);
                s10(54) <= s9(60);
                s10(55) <= s9(61);
                s10(56) <= s9(10);
                s10(57) <= s9(12);
                s10(58) <= s9(14);
                s10(59) <= s9(15);
                s10(60) <= s9(26);
                s10(61) <= s9(28);
                s10(62) <= s9(30);
                s10(63) <= s9(31);
                s10(64) <= s9(35);
                s10(65) <= s9(37);
                s10(66) <= s9(40);
                s10(67) <= s9(42);
                s10(68) <= s9(78);
                s10(69) <= s9(79);
                s10(70) <= s9(55);
                s10(71) <= s9(56);
                s10(72) <= s9(58);
                s10(73) <= s9(59);
                s11(0) <= 0.35355339059 * s10(0);
                s11(1) <= 0.35355339059 * s10(5);
                s11(2) <= 0.35355339059 * s10(6);
                s11(3) <= s10(56) + s10(7);
                s11(4) <= s10(57) + s10(8);
                s11(5) <= s10(58) + s10(7);
                s11(6) <= s10(59) + s10(8);
                s11(7) <= s10(9) + s10(10);
                s11(8) <= s10(11) + s10(12);
                s11(9) <= s10(13) + s10(14);
                s11(10) <= s10(15) + s10(16);
                s11(11) <= 0.35355339059 * s10(17);
                s11(12) <= s10(18) + s10(19);
                s11(13) <= s10(20) + s10(21);
                s11(14) <= s10(22) + s10(23);
                s11(15) <= s10(24) + s10(25);
                s11(16) <= s10(60) + s10(26);
                s11(17) <= s10(61) + s10(27);
                s11(18) <= s10(62) + s10(26);
                s11(19) <= s10(63) + s10(27);
                s11(20) <= 0.54119610014 * s10(30);
                s11(21) <= s10(64) + s10(31);
                s11(22) <= s10(65) + s10(32);
                s11(23) <= s10(66) + s10(34);
                s11(24) <= s10(67) + s10(35);
                s11(25) <= 0.54119610014 * s10(37);
                s11(26) <= s10(9) - s10(10);
                s11(27) <= s10(13) - s10(14);
                s11(28) <= s10(18) - s10(19);
                s11(29) <= s10(22) - s10(23);
                s11(30) <= 0.35355339059 * s10(40);
                s11(31) <= 0.35355339059 * s10(45);
                s11(32) <= s10(11) - s10(12);
                s11(33) <= s10(15) - s10(16);
                s11(34) <= s10(20) - s10(21);
                s11(35) <= s10(24) - s10(25);
                s11(36) <= s10(70) + s10(31);
                s11(37) <= s10(71) + s10(32);
                s11(38) <= s10(72) + s10(34);
                s11(39) <= s10(73) + s10(35);
                s11(40) <= 0.35355339059 * s10(52);
                s11(41) <= 0.35355339059 * s10(53);
                s11(42) <= s10(54);
                s11(43) <= s10(1);
                s11(44) <= s10(2);
                s11(45) <= s10(55);
                s11(46) <= s10(3);
                s11(47) <= s10(4);
                s11(48) <= s10(28);
                s11(49) <= s10(29);
                s11(50) <= s10(33);
                s11(51) <= s10(36);
                s11(52) <= s10(38);
                s11(53) <= s10(39);
                s11(54) <= s10(68);
                s11(55) <= s10(41);
                s11(56) <= s10(42);
                s11(57) <= s10(69);
                s11(58) <= s10(43);
                s11(59) <= s10(44);
                s11(60) <= s10(46);
                s11(61) <= s10(47);
                s11(62) <= s10(48);
                s11(63) <= s10(49);
                s11(64) <= s10(50);
                s11(65) <= s10(51);
                s12(0) <= s11(3) + s11(4);
                s12(1) <= s11(5) + s11(6);
                s12(2) <= s11(7) + s11(8);
                s12(3) <= s11(9) + s11(10);
                s12(4) <= s11(12) + s11(13);
                s12(5) <= s11(14) + s11(15);
                s12(6) <= s11(16) + s11(17);
                s12(7) <= s11(18) + s11(19);
                s12(8) <= s11(49) + s11(20);
                s12(9) <= 0.35355339059 * s11(21);
                s12(10) <= 0.35355339059 * s11(22);
                s12(11) <= 0.35355339059 * s11(23);
                s12(12) <= 0.35355339059 * s11(24);
                s12(13) <= s11(51) + s11(25);
                s12(14) <= s11(3) - s11(4);
                s12(15) <= 0.5 * s11(26);
                s12(16) <= 0.5 * s11(27);
                s12(17) <= 0.5 * s11(28);
                s12(18) <= 0.5 * s11(29);
                s12(19) <= s11(16) - s11(17);
                s12(20) <= s11(5) - s11(6);
                s12(21) <= 0.5 * s11(32);
                s12(22) <= 0.5 * s11(33);
                s12(23) <= 0.5 * s11(34);
                s12(24) <= 0.5 * s11(35);
                s12(25) <= s11(18) - s11(19);
                s12(26) <= s11(63) + s11(20);
                s12(27) <= 0.35355339059 * s11(36);
                s12(28) <= 0.35355339059 * s11(37);
                s12(29) <= 0.35355339059 * s11(38);
                s12(30) <= 0.35355339059 * s11(39);
                s12(31) <= s11(65) + s11(25);
                s12(32) <= s11(7) - s11(8);
                s12(33) <= s11(9) - s11(10);
                s12(34) <= s11(12) - s11(13);
                s12(35) <= s11(14) - s11(15);
                s12(36) <= s11(42);
                s12(37) <= s11(0);
                s12(38) <= s11(43);
                s12(39) <= s11(44);
                s12(40) <= s11(45);
                s12(41) <= s11(46);
                s12(42) <= s11(47);
                s12(43) <= s11(1);
                s12(44) <= s11(2);
                s12(45) <= s11(11);
                s12(46) <= s11(48);
                s12(47) <= s11(50);
                s12(48) <= s11(52);
                s12(49) <= s11(53);
                s12(50) <= s11(54);
                s12(51) <= s11(30);
                s12(52) <= s11(55);
                s12(53) <= s11(56);
                s12(54) <= s11(57);
                s12(55) <= s11(58);
                s12(56) <= s11(59);
                s12(57) <= s11(31);
                s12(58) <= s11(60);
                s12(59) <= s11(61);
                s12(60) <= s11(62);
                s12(61) <= s11(64);
                s12(62) <= s11(40);
                s12(63) <= s11(41);
                s13(0) <= s12(0) + s12(1);
                s13(1) <= 0.35355339059 * s12(2);
                s13(2) <= 0.35355339059 * s12(3);
                s13(3) <= 0.35355339059 * s12(4);
                s13(4) <= 0.35355339059 * s12(5);
                s13(5) <= s12(6) + s12(7);
                s13(6) <= 0.35355339059 * s12(8);
                s13(7) <= 0.35355339059 * s12(13);
                s13(8) <= 0.5 * s12(14);
                s13(9) <= 0.5 * s12(19);
                s13(10) <= 0.5 * s12(20);
                s13(11) <= 0.5 * s12(25);
                s13(12) <= 0.35355339059 * s12(26);
                s13(13) <= 0.35355339059 * s12(31);
                s13(14) <= s12(0) - s12(1);
                s13(15) <= 0.35355339059 * s12(32);
                s13(16) <= 0.35355339059 * s12(33);
                s13(17) <= 0.35355339059 * s12(34);
                s13(18) <= 0.35355339059 * s12(35);
                s13(19) <= s12(6) - s12(7);
                s13(20) <= s12(36);
                s13(21) <= s12(37);
                s13(22) <= s12(38);
                s13(23) <= s12(39);
                s13(24) <= s12(40);
                s13(25) <= s12(41);
                s13(26) <= s12(42);
                s13(27) <= s12(43);
                s13(28) <= s12(44);
                s13(29) <= s12(45);
                s13(30) <= s12(46);
                s13(31) <= s12(9);
                s13(32) <= s12(10);
                s13(33) <= s12(47);
                s13(34) <= s12(11);
                s13(35) <= s12(12);
                s13(36) <= s12(48);
                s13(37) <= s12(15);
                s13(38) <= s12(16);
                s13(39) <= s12(49);
                s13(40) <= s12(17);
                s13(41) <= s12(18);
                s13(42) <= s12(50);
                s13(43) <= s12(51);
                s13(44) <= s12(52);
                s13(45) <= s12(53);
                s13(46) <= s12(54);
                s13(47) <= s12(55);
                s13(48) <= s12(56);
                s13(49) <= s12(57);
                s13(50) <= s12(58);
                s13(51) <= s12(21);
                s13(52) <= s12(22);
                s13(53) <= s12(59);
                s13(54) <= s12(23);
                s13(55) <= s12(24);
                s13(56) <= s12(60);
                s13(57) <= s12(27);
                s13(58) <= s12(28);
                s13(59) <= s12(61);
                s13(60) <= s12(29);
                s13(61) <= s12(30);
                s13(62) <= s12(62);
                s13(63) <= s12(63);
                s14(0) <= 0.35355339059 * s13(0);
                s14(1) <= 0.35355339059 * s13(5);
                s14(2) <= 0.35355339059 * s13(14);
                s14(3) <= 0.35355339059 * s13(19);
                s14(4) <= s13(20);
                s14(5) <= s13(21);
                s14(6) <= s13(22);
                s14(7) <= s13(23);
                s14(8) <= s13(24);
                s14(9) <= s13(25);
                s14(10) <= s13(26);
                s14(11) <= s13(27);
                s14(12) <= s13(28);
                s14(13) <= s13(1);
                s14(14) <= s13(2);
                s14(15) <= s13(29);
                s14(16) <= s13(3);
                s14(17) <= s13(4);
                s14(18) <= s13(30);
                s14(19) <= s13(6);
                s14(20) <= s13(31);
                s14(21) <= s13(32);
                s14(22) <= s13(33);
                s14(23) <= s13(34);
                s14(24) <= s13(35);
                s14(25) <= s13(7);
                s14(26) <= s13(36);
                s14(27) <= s13(8);
                s14(28) <= s13(37);
                s14(29) <= s13(38);
                s14(30) <= s13(39);
                s14(31) <= s13(40);
                s14(32) <= s13(41);
                s14(33) <= s13(9);
                s14(34) <= s13(42);
                s14(35) <= s13(43);
                s14(36) <= s13(44);
                s14(37) <= s13(45);
                s14(38) <= s13(46);
                s14(39) <= s13(47);
                s14(40) <= s13(48);
                s14(41) <= s13(49);
                s14(42) <= s13(50);
                s14(43) <= s13(10);
                s14(44) <= s13(51);
                s14(45) <= s13(52);
                s14(46) <= s13(53);
                s14(47) <= s13(54);
                s14(48) <= s13(55);
                s14(49) <= s13(11);
                s14(50) <= s13(56);
                s14(51) <= s13(12);
                s14(52) <= s13(57);
                s14(53) <= s13(58);
                s14(54) <= s13(59);
                s14(55) <= s13(60);
                s14(56) <= s13(61);
                s14(57) <= s13(13);
                s14(58) <= s13(62);
                s14(59) <= s13(15);
                s14(60) <= s13(16);
                s14(61) <= s13(63);
                s14(62) <= s13(17);
                s14(63) <= s13(18);

            end if;
        end if;
    end process;
end architecture;
