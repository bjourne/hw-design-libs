`include "full_adder.sv"
module full_adder_tb();
endmodule
